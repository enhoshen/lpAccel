package COM;
    typedef struct packed{
    
    } fiforam_in;
endpackage
