`include "/home/enhoshen/research/lpAccel/src/MEM/MEMdefine.sv"
`include "/home/enhoshen/research/lpAccel/src/MEM/MEM.sv"
`include "/home/enhoshen/research/lpAccel/src/MEM/memv/MEMV_include.sv"

