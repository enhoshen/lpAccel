package BufCfg ;
    parameter DWD =16;
    parameter GBUFDWD=32;
    parameter IBUFSIZE=512;
    parameter WBUFSIZE=256; 
    parameter IBUFBANK=16;
    parameter WBUFBANK=16;
    parameter GBUFSIZE=1024;
    parameter GBUFBANK=32;
endpackage
