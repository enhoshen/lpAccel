import PECfg::*;

module PathStageController (
);
endmodule
