import PECfg::*;

module DataPathController(



);
endmodule
