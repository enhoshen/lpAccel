
`include "../src/define.sv"
`include "../src/PE/PEdefine.sv"
//`include "../src/PE/Aunit.sv"
//`include "../src/PE/MultADTbooth.sv"
`include "../src/common/LoopCounter.sv"
`include "../src/PE/DatapathControl.sv"

