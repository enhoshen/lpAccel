module RowAddressController #(
)(
);
endmodule
