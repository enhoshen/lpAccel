`timescale 1 ns/1 ps
`include "MEM.sv"
`include "RF_2P_48x16.v"
`include "RF_2P_48x64.v"
//`include "RF_2P_12x16.v"
`include "RF_2P_12x32.v"

