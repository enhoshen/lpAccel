module FIFORAM{
input            pop
input    
};


endmodule
