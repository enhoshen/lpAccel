import PECfg::*;

module InStageController(



);
endmodule

module DataPathController(



);
endmodule
