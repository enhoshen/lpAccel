package BufCfg ;
    parameter DWD =16;
    parameter GBUFDWD=32;
    parameter IBUFSIZE=512;
    parameter WBUFSIZE=256; 
    parameter IBUFBANK=1;
    parameter WBUFBANK=1;
    parameter GBUFSIZE=800;
    parameter GBUFBANK=2;
endpackage
