module Aunit(
input AuCtl i_ctl,
input [DWD-1:0] 
input [DWD-1:0]
);

 
