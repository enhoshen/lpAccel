module ColumnAlligner #(
)(
);
endmodule
