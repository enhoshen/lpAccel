module IF_PAD #(
)(
);
endmodule


module W_PAD #(
)(
);
endmodule


module 
