import PECfg::*;
module InputBuffer #(

)(
input [DWD-1:0] i_ 
);
endmodule
