
`include "../src/define.sv"
`include "../src/common/CommonDefine.sv"
`include "../src/MEM/MEMdefine.sv"
`include "../src/PE/PEdefine.sv"
`include "../src/common/LoopCounter.sv"
`include "../src/common/Controllers.sv"
`include "../src/PE/DatapathControl.sv"
