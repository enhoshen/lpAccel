module XBunit#(
parameter BW_O=3
parameter BW_I= 
)(
input []
input []
input []
input i_bc_se
output [] o_out 
);

logic [] xnor;
logic [] x_and;
logic [] bit_count;

assign o_out = bit_count

endmodule



