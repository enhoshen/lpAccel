module PriorityRoundRobin #(
parameter N = 3
)(
input
output 
);
endmodule

