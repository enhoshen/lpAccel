`include `"`HOME/syn/`GATE_LEVEL`"
module `GATE_LEVEL;

`TESTMODULE dut();

`default_Nico_init_block(`GATE_LEVEL,10000);
endmodule
