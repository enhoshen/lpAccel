import PECfg::*;

module PathStage(
);
endmodule
