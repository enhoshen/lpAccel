`include "../src/define.sv"
`include "../src/PE/PEdefine.sv"
`include "../src/PE/Aunit.sv"
