`include "MEMdefine.sv"
`include "MEM.sv"
`include "MEMV_include.sv"

