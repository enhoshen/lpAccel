`include "../src/define.sv"
`include "../src/PE/PEdefine.sv"
`include "../src/common/LoopCtrl.sv"
