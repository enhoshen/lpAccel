`include "../src/PE/PE_include.sv"
`include "../src/typedef.sv"
`include "../src/IF/IF.sv"
