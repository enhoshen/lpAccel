module WeightBuffer #(
)(
);
endmodule
