package COMM;
    
    function overflow 
        input a;
        begin
        end
    endfunction
    typedef struct packed{
        logic   pop,
        logic   write
    } fiforam_in;
    
endpackage
